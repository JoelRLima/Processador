LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY ROM IS
PORT(
           clock : IN STD_LOGIC; 
           rom_enable : IN STD_LOGIC;
           address : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- mudar para 15 downto 0?
           data_output : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
);
END ROM;
ARCHITECTURE behav OF ROM IS
     TYPE rom_type IS ARRAY(0 to 16) OF STD_LOGIC_VECTOR(15 DOWNTO 0); -- 16 endereços de 16 bits (utilizar 15 downto 0?)
	  
    --- INSTRUÇÕES
    --- CARREGAR: 0000 R3R2R1R0 D7D6D5D4D3D2D1D0 
    --- ARMAZENAR: 0001 R3R2R1R0 D7D6D5D4D3D2D1D0
    --- SOMAR: 0010 RA3RA2RA1RA0 RB3RB2RB1RB0 RC3RC2RC1RC0
    --- CARREGAR CONSTANTE: 0011 R3R2R1R0 C7C6C5C4C3C2C1C0
    --- SUBTRAIR: 0100 RA3RA2RA1RA0 RB3RB2RB1RB0 RC3RC2RC1RC0
    --- SALTAR SE ZERO: 0101 RA3RA2RA1RA0 O7O6O5O4O3O2O1O0
	 --- ANDbitabit: 0110 RA3RA2RA1RA0 RB3RB2RB1RB0 RC3RC2RC1RC0 ESCREVE NO RC
	 --- ORbitabit: 0111 RA3RA2RA1RA0 RB3RB2RB1RB0 RC3RC2RC1RC0 ESCREVE NO RC
	 --- NOT A: 1000 "Dont care" RB3RB2RB1RB0 RC3RC2RC1RC0 ESCREVE NO RC
     CONSTANT mem: rom_type := (
        0 => "0011000100000011", -- RF[0001]=00000011 					-- RF[0001]=3
        1 => "0011001000000010", -- RF[0010]=00000010 					-- RF[0010]=2
        2 => "0010001100010010", -- RF[0011]=RF[0001]+RF[0010] 		-- RF[0011]=3+2=5
        3 => "0001001100000001", -- D[00000001]=RF[0011]					-- D[00000001]=RF[0011]=5
		  4 => "0110001100010000", -- RF[0000]=RF[0011] AND RF[0001] 	-- RF[0000]=101 AND 011 = 001
		  5 => "0001000000000001", -- D[00000001]=RF[0000]					-- D[00000001]=001
		  6 => "0000001000000001", -- RF[0010]=D[00000001]					-- RF[0010]=001
		  7 => "0001001000000010", -- D[00000010]=RF[0010]					-- D[00000010]=001
		  8 => "0101001000000011", -- IF RF[0010]=0 THEN jump 3 positions -- 001 != 000 entao nao pula
		  9 => "0111001000110001", -- RF[0001]=RF[0010] OR RF[0011]		-- RF[0001]=001 OR 101 = 101
		  10=> "0001000100000000", -- D[00000000]=RF[0001]					-- D[00000000]=101
		  11=> "1000000000010000", -- RF[0000]= NOT(RF[0001])				-- RF[0000]= not(101)
		  12=> "0001000000000001", -- D[00000001]=RF[0000]					-- D[00000001]="1111111111111010"
		  13=> "0011001100000011", -- Load 3 into RF[0011]
		  14=> "0011000100000010", -- Load 2 into RF[0001]
		  15=> "0100000000110001", -- RF[0000]=RF[0011]-RF[0001]
		  16=> "0001000000000000", -- D[00000000]=RF[0000]
        others => "0000000000000000"
            );

BEGIN

PROCESS(clock) IS
BEGIN
    IF (RISING_EDGE(clock) AND rom_enable = '1') THEN
            data_output <= mem(conv_integer(unsigned(address)));
    END IF;
END PROCESS;
END behav;
